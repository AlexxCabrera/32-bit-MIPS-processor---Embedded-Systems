/*INCOMPLETE*/
//Dont know size for address, write data, or Read data
module DataMem(input MemWrite, MemRead, Address, Write_data
output Read_data );


endmodule
