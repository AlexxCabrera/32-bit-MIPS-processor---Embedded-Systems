/*taking ones compliment if sub is high.
This is the only way I knew how to do it.
*/
module thirtytwoBitXOR(
input	[31:0] B, [0:0] Sub,
output	[31:0] Out);

assign Out[0] = B[0] ^ Sub;
assign Out[1] = B[1] ^ Sub;
assign Out[2] = B[2] ^ Sub;
assign Out[3] = B[3] ^ Sub;
assign Out[4] = B[4] ^ Sub;
assign Out[5] = B[5] ^ Sub;
assign Out[6] = B[6] ^ Sub;
assign Out[7] = B[7] ^ Sub;
assign Out[8] = B[8] ^ Sub;
assign Out[9] = B[9] ^ Sub;
assign Out[10] = B[10] ^ Sub;
assign Out[11] = B[11] ^ Sub;
assign Out[12] = B[12] ^ Sub;
assign Out[13] = B[13] ^ Sub;
assign Out[14] = B[14] ^ Sub;
assign Out[15] = B[15] ^ Sub;
assign Out[16] = B[16] ^ Sub;
assign Out[17] = B[17] ^ Sub;
assign Out[18] = B[18] ^ Sub;
assign Out[19] = B[19] ^ Sub;
assign Out[20] = B[20] ^ Sub;
assign Out[21] = B[21] ^ Sub;
assign Out[22] = B[22] ^ Sub;
assign Out[23] = B[23] ^ Sub;
assign Out[24] = B[24] ^ Sub;
assign Out[25] = B[25] ^ Sub;
assign Out[26] = B[26] ^ Sub;
assign Out[27] = B[27] ^ Sub;
assign Out[28] = B[28] ^ Sub;
assign Out[29] = B[29] ^ Sub;
assign Out[30] = B[30] ^ Sub;
assign Out[31] = B[31] ^ Sub;
	
endmodule
