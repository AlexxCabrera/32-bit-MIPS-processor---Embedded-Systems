/*32-BITWISE OR*/
module Or_32 (Y, A, B);
input [31:0] A, B;
output [31:0] Y;

	Or o0(.Y(Y[0]),.A(A[0]),.B(B[0]));
	Or o1(.Y(Y[1]),.A(A[1]),.B(B[1]));
	Or o2(.Y(Y[2]),.A(A[2]),.B(B[2]));
	Or o3(.Y(Y[3]),.A(A[3]),.B(B[3]));
	Or o4(.Y(Y[4]),.A(A[4]),.B(B[4]));
	Or o5(.Y(Y[5]),.A(A[5]),.B(B[5]));
	Or o6(.Y(Y[6]),.A(A[6]),.B(B[6]));
	Or o7(.Y(Y[7]),.A(A[7]),.B(B[7]));
	Or o8(.Y(Y[8]),.A(A[8]),.B(B[8]));
	Or o9(.Y(Y[9]),.A(A[9]),.B(B[9]));
	Or o10(.Y(Y[10]),.A(A[10]),.B(B[10]));
	Or o11(.Y(Y[11]),.A(A[11]),.B(B[11]));
	Or o12(.Y(Y[12]),.A(A[12]),.B(B[12]));
	Or o13(.Y(Y[13]),.A(A[13]),.B(B[13]));
	Or o14(.Y(Y[14]),.A(A[14]),.B(B[14]));
	Or o15(.Y(Y[15]),.A(A[15]),.B(B[15]));
	Or o16(.Y(Y[16]),.A(A[16]),.B(B[16]));
	Or o17(.Y(Y[17]),.A(A[17]),.B(B[17]));
	Or o18(.Y(Y[18]),.A(A[18]),.B(B[18]));
	Or o19(.Y(Y[19]),.A(A[19]),.B(B[19]));
	Or o20(.Y(Y[20]),.A(A[20]),.B(B[20]));
	Or o21(.Y(Y[21]),.A(A[21]),.B(B[21]));
	Or o22(.Y(Y[22]),.A(A[22]),.B(B[22]));
	Or o23(.Y(Y[23]),.A(A[23]),.B(B[23]));
	Or o24(.Y(Y[24]),.A(A[24]),.B(B[24]));
	Or o25(.Y(Y[25]),.A(A[25]),.B(B[25]));
	Or o26(.Y(Y[26]),.A(A[26]),.B(B[26]));
	Or o27(.Y(Y[27]),.A(A[27]),.B(B[27]));
	Or o28(.Y(Y[28]),.A(A[28]),.B(B[28]));
	Or o29(.Y(Y[29]),.A(A[29]),.B(B[29]));
	Or o30(.Y(Y[30]),.A(A[30]),.B(B[30]));
	Or o31(.Y(Y[31]),.A(A[31]),.B(B[31]));

endmodule 
