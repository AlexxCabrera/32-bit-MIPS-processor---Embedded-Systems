module ShiftLeft2(output out, input [31:0] in);

assign out = in<<2;

endmodule 
