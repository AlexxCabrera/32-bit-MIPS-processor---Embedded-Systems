module Instruction_memory(input ReadAddress, output	[31:0] instruction);


	
endmodule 
