/*INCOMPLETE*/
module Instruction_memory(input [31:0] ReadAddress, output[31:0] instruction);


	
endmodule 
