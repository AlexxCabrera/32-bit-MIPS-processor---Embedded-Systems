/*INCOMPLETE*/
module Control(input [5:0] instruction, output RegDst, Branch, MemRead, MemtoReg,ALUOp, MemWrite, ALUSrc, RegWrite);
	
endmodule 
