module or_32tb;
	wire [31:0] Y;
	reg [31:0] A, B;

	Or_32 or32_tb(Y,A,B);

	initial begin
		A = 32'b00010111111100010011111011101000;	B = 32'b10110000100110010111111100000111;	#5; //10110111111110010111111111101111
		A = 32'b00000000000000000000000000000000;	B = 32'b10110000100110010111111100000111;	#5; //10110000100110010111111100000111
		A = 32'b11111111111111111111111111111111;	B = 32'b10110000100110010111111100000111;	#5; //11111111111111111111111111111111
		A = 32'b01010001001110110001000001010010;	B = 32'b00001111111100011100111000100101;	#5; //01011111111110111101111001110111
	end

	initial begin
		$monitor("Y = %b",Y);
	end


endmodule
