/*INCOMPLETE*/
module RegDstMux(input clk, [4:0] read_register1, [4:0] read_register2, [4:0] writeReg, [0:0] RegWrite, [31:0] writeData, 
output reg [31:0] readData1, readData2);

reg [31:0] registers [31:0];

endmodule
